module Mem(clock, dataWB_enable, dataWB_data);

input clock, dataWB_enable;
input[16:0] dataWB_data;
reg[16:0]data[3:0];

//StateMachine st0
//StateMachine st1
//StateMachine st2
//StateMachine st3


endmodule
