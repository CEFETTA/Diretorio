module Diretorio (clock);

Mem M0(clock, dataWB_enable, dataWB_data);




endmodule
